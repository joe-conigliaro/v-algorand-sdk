module crypto2

const (
	err_invalid_signature_returned         = error('ed25519 library returned an invalid signature')
	err_invalid_private_key                = error('invalid private key')
	err_msig_unknown_version               = error('unknown version != 1')
	err_msig_invalid_threshold             = error('invalid threshold')
	err_msig_invalid_secret_key            = error('secret key has no corresponding public identity in multisig preimage')
	err_msig_merge_less_than_two           = error('cannot merge fewer than two multisig transactions')
	err_msig_merge_keys_mismatch           = error('multisig parameters do not match')
	err_msig_merge_invalid_dups            = error('mismatched duplicate signatures')
	err_msig_merge_auth_addr_mismatch      = error('mismatched AuthAddrs')
	err_lsig_too_many_signatures           = error('logicsig has too many signatures, at most one of Sig or Msig may be defined')
	err_lsig_no_signature                  = error('logicsig is not delegated')
	err_lsig_invalid_signature             = error('invalid logicsig signature')
	err_lsig_no_public_key                 = error('missing public key of delegated logicsig')
	err_lsig_invalid_public_key            = error('public key does not match logicsig signature')
	err_lsig_invalid_program               = error('invalid logicsig program')
	err_lsig_empty_msig                    = error('empty multisig in logicsig')
	err_lsig_account_public_key_not_needed = error('a public key for the signer was provided when none was expected')
)
